module top_module(output one,zero);
    assign one = 0;
endmodule