module top_module (
    input d, 
    input ena,
    output q);

endmodule